`define OPCODE_ANDREG 11'b?0001010???
`define OPCODE_ORRREG 11'b?0101010???
`define OPCODE_ADDREG 11'b?0?01011???
`define OPCODE_SUBREG 11'b?1?01011???

`define OPCODE_ADDIMM 11'b?0?10001???
`define OPCODE_SUBIMM 11'b?1?10001???

`define OPCODE_MOVZ   11'b110100101??

`define OPCODE_B      11'b?00101?????
`define OPCODE_CBZ    11'b?011010????

`define OPCODE_LDUR   11'b??111000010
`define OPCODE_STUR   11'b??111000000

module control(
	       output reg 	reg2loc,
	       output reg 	alusrc,
	       output reg 	mem2reg,
	       output reg 	regwrite,
	       output reg 	memread,
	       output reg 	memwrite,
	       output reg 	branch,
	       output reg 	uncond_branch,
	       output reg [3:0] aluop,
	       output reg [2:0] signop, // changed to be 3 bits for MOVZ
	       input [10:0] 	opcode
	       );

   always @(*)
     begin
	casez (opcode)

          /* Add cases here for each instruction your processor supports */
	 
	  `OPCODE_LDUR: // LDUR (D instruction)
	    begin
	       reg2loc       = 1'bx;
               uncond_branch = 1'b0;
               branch        = 1'b0;
               memread       = 1'b1;
               mem2reg       = 1'b1;
               memwrite      = 1'b0;
               alusrc        = 1'b1;
               regwrite      = 1'b1;
               aluop         = 4'b0010;
               signop        = 3'b010;
               $display("LDUR received");
	    end // case: `OPCODE_LDUR

	  `OPCODE_STUR: // STUR (D instruction)
	    begin
	       reg2loc       = 1'b1;
               uncond_branch = 1'b0;
               branch        = 1'b0;
               memread       = 1'b0;
               mem2reg       = 1'bx;
               memwrite      = 1'b1;
               alusrc        = 1'b1;
               regwrite      = 1'b0;
               aluop         = 4'b0010;
               signop        = 3'b010;
               $display("STUR received");
	    end // case: `OPCODE_STUR

	  `OPCODE_ADDREG: // ADDR (R instruction)
	    begin
	       reg2loc       = 1'b0;
               uncond_branch = 1'b0;
               branch        = 1'b0;
               memread       = 1'b0;
               mem2reg       = 1'b0;
               memwrite      = 1'b0;
               alusrc        = 1'b0;
               regwrite      = 1'b1;
               aluop         = 4'b0010;
               signop        = 3'bxxx;
               $display("ADDR received");
	    end // case: `OPCODE_ADDREG

	  `OPCODE_ADDIMM: // ADDI (I instruction)
	    begin
	       reg2loc       = 1'b0;
               uncond_branch = 1'b0;
               branch        = 1'b0;
               memread       = 1'b0;
               mem2reg       = 1'b0;
               memwrite      = 1'b0;
               alusrc        = 1'b0;
               regwrite      = 1'b1;
               aluop         = 4'b0010;
               signop        = 3'b011;
               $display("ADDI received");
	    end // case: `OPCODE_ADDIMM

	  `OPCODE_SUBREG: // SUBR (R instruction)
	    begin
	       reg2loc       = 1'b0;
               uncond_branch = 1'b0;
               branch        = 1'b0;
               memread       = 1'b0;
               mem2reg       = 1'b0;
               memwrite      = 1'b0;
               alusrc        = 1'b0;
               regwrite      = 1'b1;
               aluop         = 4'b0110;
               signop        = 3'bxxx;
               $display("SUBR received");
	    end // case: `OPCODE_SUBREG

	  `OPCODE_SUBIMM: // SUBI (I instruction)
	    begin
	       
	       reg2loc       = 1'b0;
               uncond_branch = 1'b0;
               branch        = 1'b0;
               memread       = 1'b0;
               mem2reg       = 1'b0;
               memwrite      = 1'b0;
               alusrc        = 1'b0;
               regwrite      = 1'b1;
               aluop         = 4'b0110;
               signop        = 3'b011;
               $display("SUBI received");
	    end // case: `OPCODE_SUBIMM

	  `OPCODE_ANDREG: // AND (R instruction)
	    begin
	       reg2loc       = 1'b0;
               uncond_branch = 1'b0;
               branch        = 1'b0;
               memread       = 1'b0;
               mem2reg       = 1'b0;
               memwrite      = 1'b0;
               alusrc        = 1'b0;
               regwrite      = 1'b1;
               aluop         = 4'b0000;
               signop        = 3'bxxx;
               $display("AND received");
	    end // case: `OPCODE_ANDREG

	  `OPCODE_ORRREG: // ORR (R instruction)
	    begin
	       reg2loc       = 1'b0;
               uncond_branch = 1'b0;
               branch        = 1'b0;
               memread       = 1'b0;
               mem2reg       = 1'b0;
               memwrite      = 1'b0;
               alusrc        = 1'b0;
               regwrite      = 1'b1;
               aluop         = 4'b0001;
               signop        = 3'bxxx;
               $display("ORR received");
	    end // case: `OPCODE_ORRREG

	  `OPCODE_CBZ: // CBZ (CBZ instruction)
	    begin
	       reg2loc       = 1'b1;
               uncond_branch = 1'b0;
               branch        = 1'b1;
               memread       = 1'b0;
               mem2reg       = 1'bx;
               memwrite      = 1'b0;
               alusrc        = 1'b0;
               regwrite      = 1'b0;
               aluop         = 4'b0111;
               signop        = 3'b001;
               $display("CBZ received");
	    end // case: `OPCODE_CBZ

	  `OPCODE_B: // B (B instruction)
	    begin
	       reg2loc       = 1'bx;
               uncond_branch = 1'b1;
               branch        = 1'bx;
               memread       = 1'b0;
               mem2reg       = 1'bx;
               memwrite      = 1'b0;
               alusrc        = 1'bx;
               regwrite      = 1'b0;
               aluop         = 4'bxxxx;
               signop        = 3'b000;
               $display("B received");
	    end // case: `OPCODE_B

	  `OPCODE_MOVZ: // MOVZ 1 (IM instruction)
	    begin
	       // IMPLEMENT:
	       reg2loc       = 1'bx;
               uncond_branch = 1'b0;
               branch        = 1'b0;
               memread       = 1'b0;
               mem2reg       = 1'b0;
               memwrite      = 1'b0;
               alusrc        = 1'b1;
               regwrite      = 1'b1;
               aluop         = 4'b0111;
               signop        = opcode[2:0]; //opcode[2:0]
               $display("MOVZ received");
	    end // case: `OPCODE_MOVZ
       
	endcase // casez (opcode)
	
     end // always @ (*)
endmodule

